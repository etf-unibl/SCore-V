-----------------------------------------------------------------------------
-- Faculty of Electrical Engineering
-- PDS 2025
-- https://github.com/etf-unibl/pds-2025/
-----------------------------------------------------------------------------
--
-- unit name:     pc_next_instruction
--
-- description:
--
--   This file implements a simple next Program Counter (PC) calculation
--   logic.
--
-----------------------------------------------------------------------------
-- Copyright (c) 2025 Faculty of Electrical Engineering
-----------------------------------------------------------------------------
-- The MIT License
-----------------------------------------------------------------------------
-- Copyright 2025 Faculty of Electrical Engineering
--
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the "Software"),
-- to deal in the Software without restriction, including without limitation
-- the rights to use, copy, modify, merge, publish, distribute, sublicense,
-- and/or sell copies of the Software, and to permit persons to whom
-- the Software is furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
-- THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,
-- ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
-- OTHER DEALINGS IN THE SOFTWARE
-----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--! @file pc_next_instruction.vhd
--! @brief Next sequential Program Counter calculation
--! @details Computes the next instruction address by incrementing
--! the current PC value by 4.

entity pc_next_instruction is
  port (
    pc_i       : in  std_logic_vector(31 downto 0); --! Current Program Counter value
    pc_next_o  : out std_logic_vector(31 downto 0)  --! Next sequential PC value
  );
end pc_next_instruction;

--! @brief Architecture arch for next PC computation
--! @details Implements combinational logic for sequential PC increment.
architecture arch of pc_next_instruction is
  --! @brief Internal signal declarations
  signal tmp : unsigned(31 downto 0); --! Temporary unsigned signal for arithmetic operation
begin
  tmp <= unsigned(pc_i) + 4;
  
  --! @brief Output assignment
  pc_next_o <= std_logic_vector(tmp);
end arch;
