-----------------------------------------------------------------------------
-- Faculty of Electrical Engineering
-- PDS 2025
-- https://github.com/etf-unibl/SCore-V
-----------------------------------------------------------------------------
--
-- unit name:     counter_vunit_example
--
-- description:
--
--   This file implements a simple counter used for showcasing VUnit test
--
-----------------------------------------------------------------------------
-- Copyright (c) 2025 Faculty of Electrical Engineering
-----------------------------------------------------------------------------
-- The MIT License
-----------------------------------------------------------------------------
-- Copyright 2025 Faculty of Electrical Engineering
--
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the "Software"),
-- to deal in the Software without restriction, including without limitation
-- the rights to use, copy, modify, merge, publish, distribute, sublicense,
-- and/or sell copies of the Software, and to permit persons to whom
-- the Software is furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
-- THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,
-- ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
-- OTHER DEALINGS IN THE SOFTWARE
-----------------------------------------------------------------------------

-----------------------------------------------------------------------------
--! @file counter_vunit_example.vhd
--! @brief Implements a simple counter used to demonstrate vunit tests
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--! @brief Entity definition of counter_vunit_example
--! Unit implements a simple 4-bit counter.
entity counter_vunit_example is
  port (
    clk_i    : in  std_logic;                   --! Clock input of the unit
    rst_i    : in  std_logic;                   --! Reset input of the unit
    enable_i : in  std_logic;                   --! Input which enables counting
    count_o  : out std_logic_vector(3 downto 0) --! 4-bit output of the counter
  );
end entity counter_vunit_example;

--! @brief Architecture definition of counter_vunit_example
--! On every positive edge of clock counter increases
--! count_o by one.
architecture arch of counter_vunit_example is
  signal count_reg : unsigned(3 downto 0);
begin

  -- process main
  main : process(clk_i, rst_i)
  begin
    if rst_i = '1' then
      count_reg <= (others => '0');
    elsif rising_edge(clk_i) then
      if enable_i = '1' then
        count_reg <= count_reg + 1;
      end if;
    end if;
  end process main;

  count_o <= std_logic_vector(count_reg);

end architecture arch;
